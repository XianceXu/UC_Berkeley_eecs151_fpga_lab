// module adder()
// input 